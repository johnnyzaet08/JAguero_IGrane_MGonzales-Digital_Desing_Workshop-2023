module display_game_over(
	input wire [9:0] counter_x,
	input wire [9:0] counter_y,
	output reg [7:0] r_red,
	output reg [7:0] r_green,
	output reg [7:0] r_blue  
);

	/* Design "¡Has perdido!" message to display. The same way vga controller is programmed */

endmodule