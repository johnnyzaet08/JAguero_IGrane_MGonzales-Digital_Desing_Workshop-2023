module display_game_over(
	output wire [7:0] red_d,	    //red vga output
   output wire [7:0] green_d,     //green vga output
   output wire [7:0] blue_d	    //blue vga output
);

	/* Design "¡Has perdido!" message to display. The same way vga controller is programmed */

endmodule