`timescale 1 ns / 1 ps

module Shifting_TB();
	
	reg [3:0] a;
	wire [3:0] y;
	
	Shifting dut(a, 1, y);

	initial begin
		a = 4'b0000; #20; //0
		a = 4'b0001; #20; //1
		a = 4'b0010; #20; //2
		a = 4'b0011; #20; //3
		a = 4'b0100; #20; //4
		a = 4'b0101; #20; //5
		a = 4'b0110; #20; //6
		a = 4'b0111; #20; //7
		a = 4'b1000; #20; //8
		a = 4'b1001; #20; //0
		a = 4'b1010; #20; //10
		a = 4'b1011; #20; //11
		a = 4'b1100; #20; //12
		a = 4'b1101; #20; //13
		a = 4'b1110; #20; //14
		a = 4'b1111; #20; //15
	end

endmodule